module ajuste (r, s, y);
	input [59:0] r;
	input [5:0] s;
	output reg [17:0] y;
	
		always@(r)
		case(s)
			0 : y = r[17:0]; 
			1 : y = r[18:1]; 
			2 : y = r[19:2]; 
			3 : y = r[20:3];
			4 : y = r[21:4];
			5 :	y = r[22:5];
			6 :	y = r[23:6];
			7 : y = r[24:7];
			8 :	y = r[25:8];
			9 :	y = r[26:9];
			10 : y = r[27:10];
			11 : y = r[28:11];
			12 : y = r[29:12];
			13 : y = r[30:13];
			14 : y = r[31:14];
			15 : y = r[32:15];
			16 : y = r[33:16];
			17 : y = r[34:17];
			18 : y = r[35:18];
			19 : y = r[36:19];
			20 : y = r[37:20];
			21 : y = r[38:21];
			22 : y = r[39:22];
			23 : y = r[40:23];
			24 : y = r[41:24];
			25 : y = r[42:25];
			26 : y = r[43:26];
			27 : y = r[44:27];
			28 : y = r[45:28];
			29 : y = r[46:29];
			30 : y = r[47:30];
			31 : y = r[48:31];
			32 : y = r[49:32];
			33 : y = r[50:33];
			34 : y = r[51:34];
			35 : y = r[52:35];
			36 : y = r[53:36];
			37 : y = r[54:37];
			38 : y = r[55:38];
			39 : y = r[56:39];
			40 : y = r[57:40];
			41 : y = r[58:41];
			42 : y = r[59:42]; 
			default y = 0;
		endcase
		
endmodule